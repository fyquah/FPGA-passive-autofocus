// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: lpm_mux3.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module lpm_mux3 (
	data0x,
	data1x,
	sel,
	result);

	input	[89:0]  data0x;
	input	[89:0]  data1x;
	input	  sel;
	output	[89:0]  result;

	wire [89:0] sub_wire0;
	wire [89:0] sub_wire3 = data1x[89:0];
	wire [89:0] result = sub_wire0[89:0];
	wire [89:0] sub_wire1 = data0x[89:0];
	wire [179:0] sub_wire2 = {sub_wire3, sub_wire1};
	wire  sub_wire4 = sel;
	wire  sub_wire5 = sub_wire4;

	lpm_mux	LPM_MUX_component (
				.data (sub_wire2),
				.sel (sub_wire5),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		LPM_MUX_component.lpm_size = 2,
		LPM_MUX_component.lpm_type = "LPM_MUX",
		LPM_MUX_component.lpm_width = 90,
		LPM_MUX_component.lpm_widths = 1;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "2"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "90"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "1"
// Retrieval info: USED_PORT: data0x 0 0 90 0 INPUT NODEFVAL "data0x[89..0]"
// Retrieval info: USED_PORT: data1x 0 0 90 0 INPUT NODEFVAL "data1x[89..0]"
// Retrieval info: USED_PORT: result 0 0 90 0 OUTPUT NODEFVAL "result[89..0]"
// Retrieval info: USED_PORT: sel 0 0 0 0 INPUT NODEFVAL "sel"
// Retrieval info: CONNECT: @data 0 0 90 0 data0x 0 0 90 0
// Retrieval info: CONNECT: @data 0 0 90 90 data1x 0 0 90 0
// Retrieval info: CONNECT: @sel 0 0 1 0 sel 0 0 0 0
// Retrieval info: CONNECT: result 0 0 90 0 @result 0 0 90 0
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux3.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux3.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux3.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux3.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux3_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux3_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
